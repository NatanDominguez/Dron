



module pwm_gen #(
    parameter int BASE = 1000  
) (
    input logic clk_i,
    input logic rst_ni,

    output logic pwm_o
);



endmodule